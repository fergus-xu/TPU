module fpAdder32(
	input logic [31:0] A,
	input logic [31:0] B,
	output logic [31:0] out
);
	output [7:0] diff;
	logic EA_lt_EB;
	exponent_difference ed (A[30:23], B[30:23], )



endmodule 